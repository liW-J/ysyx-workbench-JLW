module shifter(
    input                   [31 : 0]        src0,
    input                   [ 4 : 0]        src1,
    output                  [31 : 0]        res1,       //逻辑右移
    output                  [31 : 0]        res2        //算术右移
);
// Write your code here

// End of your code
endmodule
